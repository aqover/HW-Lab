
///
/// created by p8051Rom.exe
/// author: Simon Teran (simont@opencores.org)
///
/// source file: D:\verilog\oc8051\test\sqroot.hex
/// date: 6.6.02
/// time: 22:01:15
///

module oc8051_rom (rst, clk, addr, ea_int, data1, data2, data3);

parameter INT_ROM_WID= 11;

input rst, clk;
input [15:0] addr;
output ea_int;
output [7:0] data1, data2, data3;
reg [7:0] data1, data2, data3;
reg [7:0] buff [65535:0];
integer i;

wire ea;

assign ea = | addr[15:INT_ROM_WID];
assign ea_int = ! ea;

initial
begin
    for (i=0; i<65536; i=i+1)
      buff [i] = 8'h00;
#2

    buff [16'h00_00] = 8'h02;
    buff [16'h00_01] = 8'h04;
    buff [16'h00_02] = 8'h54;
    buff [16'h00_03] = 8'h7F;
    buff [16'h00_04] = 8'h00;
    buff [16'h00_05] = 8'h7E;
    buff [16'h00_06] = 8'h00;
    buff [16'h00_07] = 8'h7D;
    buff [16'h00_08] = 8'h40;
    buff [16'h00_09] = 8'h7C;
    buff [16'h00_0a] = 8'h40;
    buff [16'h00_0b] = 8'h75;
    buff [16'h00_0c] = 8'h0B;
    buff [16'h00_0d] = 8'h00;
    buff [16'h00_0e] = 8'h75;
    buff [16'h00_0f] = 8'h0A;
    buff [16'h00_10] = 8'h00;
    buff [16'h00_11] = 8'h75;
    buff [16'h00_12] = 8'h09;
    buff [16'h00_13] = 8'h80;
    buff [16'h00_14] = 8'h75;
    buff [16'h00_15] = 8'h08;
    buff [16'h00_16] = 8'h40;
    buff [16'h00_17] = 8'hA8;
    buff [16'h00_18] = 8'h04;
    buff [16'h00_19] = 8'hA9;
    buff [16'h00_1a] = 8'h05;
    buff [16'h00_1b] = 8'hAA;
    buff [16'h00_1c] = 8'h06;
    buff [16'h00_1d] = 8'hAB;
    buff [16'h00_1e] = 8'h07;
    buff [16'h00_1f] = 8'h12;
    buff [16'h00_20] = 8'h01;
    buff [16'h00_21] = 8'h7A;
    buff [16'h00_22] = 8'h8F;
    buff [16'h00_23] = 8'h0F;
    buff [16'h00_24] = 8'h8E;
    buff [16'h00_25] = 8'h0E;
    buff [16'h00_26] = 8'h8D;
    buff [16'h00_27] = 8'h0D;
    buff [16'h00_28] = 8'h8C;
    buff [16'h00_29] = 8'h0C;
    buff [16'h00_2a] = 8'h12;
    buff [16'h00_2b] = 8'h02;
    buff [16'h00_2c] = 8'h80;
    buff [16'h00_2d] = 8'h8F;
    buff [16'h00_2e] = 8'h80;
    buff [16'h00_2f] = 8'hAF;
    buff [16'h00_30] = 8'h0B;
    buff [16'h00_31] = 8'hAE;
    buff [16'h00_32] = 8'h0A;
    buff [16'h00_33] = 8'hAD;
    buff [16'h00_34] = 8'h09;
    buff [16'h00_35] = 8'hAC;
    buff [16'h00_36] = 8'h08;
    buff [16'h00_37] = 8'hA8;
    buff [16'h00_38] = 8'h04;
    buff [16'h00_39] = 8'hA9;
    buff [16'h00_3a] = 8'h05;
    buff [16'h00_3b] = 8'hAA;
    buff [16'h00_3c] = 8'h06;
    buff [16'h00_3d] = 8'hAB;
    buff [16'h00_3e] = 8'h07;
    buff [16'h00_3f] = 8'h12;
    buff [16'h00_40] = 8'h01;
    buff [16'h00_41] = 8'h7A;
    buff [16'h00_42] = 8'h8F;
    buff [16'h00_43] = 8'h13;
    buff [16'h00_44] = 8'h8E;
    buff [16'h00_45] = 8'h12;
    buff [16'h00_46] = 8'h8D;
    buff [16'h00_47] = 8'h11;
    buff [16'h00_48] = 8'h8C;
    buff [16'h00_49] = 8'h10;
    buff [16'h00_4a] = 8'h12;
    buff [16'h00_4b] = 8'h02;
    buff [16'h00_4c] = 8'h80;
    buff [16'h00_4d] = 8'h8F;
    buff [16'h00_4e] = 8'h90;
    buff [16'h00_4f] = 8'hAF;
    buff [16'h00_50] = 8'h13;
    buff [16'h00_51] = 8'hAE;
    buff [16'h00_52] = 8'h12;
    buff [16'h00_53] = 8'hAD;
    buff [16'h00_54] = 8'h11;
    buff [16'h00_55] = 8'hAC;
    buff [16'h00_56] = 8'h10;
    buff [16'h00_57] = 8'hAB;
    buff [16'h00_58] = 8'h0F;
    buff [16'h00_59] = 8'hAA;
    buff [16'h00_5a] = 8'h0E;
    buff [16'h00_5b] = 8'hA9;
    buff [16'h00_5c] = 8'h0D;
    buff [16'h00_5d] = 8'hA8;
    buff [16'h00_5e] = 8'h0C;
    buff [16'h00_5f] = 8'h12;
    buff [16'h00_60] = 8'h00;
    buff [16'h00_61] = 8'h89;
    buff [16'h00_62] = 8'h8F;
    buff [16'h00_63] = 8'h17;
    buff [16'h00_64] = 8'h8E;
    buff [16'h00_65] = 8'h16;
    buff [16'h00_66] = 8'h8D;
    buff [16'h00_67] = 8'h15;
    buff [16'h00_68] = 8'h8C;
    buff [16'h00_69] = 8'h14;
    buff [16'h00_6a] = 8'h12;
    buff [16'h00_6b] = 8'h02;
    buff [16'h00_6c] = 8'h80;
    buff [16'h00_6d] = 8'h8F;
    buff [16'h00_6e] = 8'hA0;
    buff [16'h00_6f] = 8'hAF;
    buff [16'h00_70] = 8'h17;
    buff [16'h00_71] = 8'hAE;
    buff [16'h00_72] = 8'h16;
    buff [16'h00_73] = 8'hAD;
    buff [16'h00_74] = 8'h15;
    buff [16'h00_75] = 8'hAC;
    buff [16'h00_76] = 8'h14;
    buff [16'h00_77] = 8'h12;
    buff [16'h00_78] = 8'h03;
    buff [16'h00_79] = 8'hAE;
    buff [16'h00_7a] = 8'h12;
    buff [16'h00_7b] = 8'h02;
    buff [16'h00_7c] = 8'h80;
    buff [16'h00_7d] = 8'h8F;
    buff [16'h00_7e] = 8'hB0;
    buff [16'h00_7f] = 8'h80;
    buff [16'h00_80] = 8'hFE;
    buff [16'h00_81] = 8'h22;
    buff [16'h00_82] = 8'h02;
    buff [16'h00_83] = 8'h02;
    buff [16'h00_84] = 8'hEC;
    buff [16'h00_85] = 8'hE8;
    buff [16'h00_86] = 8'h64;
    buff [16'h00_87] = 8'h80;
    buff [16'h00_88] = 8'hF8;
    buff [16'h00_89] = 8'hE9;
    buff [16'h00_8a] = 8'h33;
    buff [16'h00_8b] = 8'hE8;
    buff [16'h00_8c] = 8'h33;
    buff [16'h00_8d] = 8'h60;
    buff [16'h00_8e] = 8'h11;
    buff [16'h00_8f] = 8'h04;
    buff [16'h00_90] = 8'h60;
    buff [16'h00_91] = 8'hF0;
    buff [16'h00_92] = 8'hED;
    buff [16'h00_93] = 8'h33;
    buff [16'h00_94] = 8'hEC;
    buff [16'h00_95] = 8'h33;
    buff [16'h00_96] = 8'h70;
    buff [16'h00_97] = 8'h09;
    buff [16'h00_98] = 8'hE8;
    buff [16'h00_99] = 8'hFC;
    buff [16'h00_9a] = 8'hE9;
    buff [16'h00_9b] = 8'hFD;
    buff [16'h00_9c] = 8'hEA;
    buff [16'h00_9d] = 8'hFE;
    buff [16'h00_9e] = 8'hEB;
    buff [16'h00_9f] = 8'hFF;
    buff [16'h00_a0] = 8'h22;
    buff [16'h00_a1] = 8'h04;
    buff [16'h00_a2] = 8'h60;
    buff [16'h00_a3] = 8'hDE;
    buff [16'h00_a4] = 8'hD3;
    buff [16'h00_a5] = 8'hEB;
    buff [16'h00_a6] = 8'h9F;
    buff [16'h00_a7] = 8'hEA;
    buff [16'h00_a8] = 8'h9E;
    buff [16'h00_a9] = 8'hE9;
    buff [16'h00_aa] = 8'h9D;
    buff [16'h00_ab] = 8'hE8;
    buff [16'h00_ac] = 8'hC2;
    buff [16'h00_ad] = 8'hE7;
    buff [16'h00_ae] = 8'h8C;
    buff [16'h00_af] = 8'hF0;
    buff [16'h00_b0] = 8'hC2;
    buff [16'h00_b1] = 8'hF7;
    buff [16'h00_b2] = 8'h95;
    buff [16'h00_b3] = 8'hF0;
    buff [16'h00_b4] = 8'h40;
    buff [16'h00_b5] = 8'h0C;
    buff [16'h00_b6] = 8'hE8;
    buff [16'h00_b7] = 8'hCC;
    buff [16'h00_b8] = 8'hF8;
    buff [16'h00_b9] = 8'hE9;
    buff [16'h00_ba] = 8'hCD;
    buff [16'h00_bb] = 8'hF9;
    buff [16'h00_bc] = 8'hEA;
    buff [16'h00_bd] = 8'hCE;
    buff [16'h00_be] = 8'hFA;
    buff [16'h00_bf] = 8'hEB;
    buff [16'h00_c0] = 8'hCF;
    buff [16'h00_c1] = 8'hFB;
    buff [16'h00_c2] = 8'h12;
    buff [16'h00_c3] = 8'h02;
    buff [16'h00_c4] = 8'hB7;
    buff [16'h00_c5] = 8'h85;
    buff [16'h00_c6] = 8'hD0;
    buff [16'h00_c7] = 8'hF0;
    buff [16'h00_c8] = 8'h58;
    buff [16'h00_c9] = 8'h04;
    buff [16'h00_ca] = 8'h70;
    buff [16'h00_cb] = 8'h03;
    buff [16'h00_cc] = 8'h20;
    buff [16'h00_cd] = 8'hD5;
    buff [16'h00_ce] = 8'hB3;
    buff [16'h00_cf] = 8'hE8;
    buff [16'h00_d0] = 8'h04;
    buff [16'h00_d1] = 8'h70;
    buff [16'h00_d2] = 8'h07;
    buff [16'h00_d3] = 8'h50;
    buff [16'h00_d4] = 8'h02;
    buff [16'h00_d5] = 8'hB2;
    buff [16'h00_d6] = 8'hD5;
    buff [16'h00_d7] = 8'h02;
    buff [16'h00_d8] = 8'h02;
    buff [16'h00_d9] = 8'hF6;
    buff [16'h00_da] = 8'h92;
    buff [16'h00_db] = 8'hD5;
    buff [16'h00_dc] = 8'hEC;
    buff [16'h00_dd] = 8'h04;
    buff [16'h00_de] = 8'h60;
    buff [16'h00_df] = 8'hF7;
    buff [16'h00_e0] = 8'hE4;
    buff [16'h00_e1] = 8'hCC;
    buff [16'h00_e2] = 8'hC0;
    buff [16'h00_e3] = 8'hE0;
    buff [16'h00_e4] = 8'hC3;
    buff [16'h00_e5] = 8'h98;
    buff [16'h00_e6] = 8'hF8;
    buff [16'h00_e7] = 8'h60;
    buff [16'h00_e8] = 8'h3B;
    buff [16'h00_e9] = 8'h94;
    buff [16'h00_ea] = 8'h18;
    buff [16'h00_eb] = 8'h60;
    buff [16'h00_ec] = 8'h08;
    buff [16'h00_ed] = 8'h40;
    buff [16'h00_ee] = 8'h0D;
    buff [16'h00_ef] = 8'hD0;
    buff [16'h00_f0] = 8'hE0;
    buff [16'h00_f1] = 8'hFB;
    buff [16'h00_f2] = 8'h02;
    buff [16'h00_f3] = 8'h02;
    buff [16'h00_f4] = 8'hCE;
    buff [16'h00_f5] = 8'hE4;
    buff [16'h00_f6] = 8'hFB;
    buff [16'h00_f7] = 8'hFA;
    buff [16'h00_f8] = 8'hC9;
    buff [16'h00_f9] = 8'hFC;
    buff [16'h00_fa] = 8'h80;
    buff [16'h00_fb] = 8'h28;
    buff [16'h00_fc] = 8'hE8;
    buff [16'h00_fd] = 8'h30;
    buff [16'h00_fe] = 8'hE4;
    buff [16'h00_ff] = 8'h06;
    buff [16'h01_00] = 8'hE4;
    buff [16'h01_01] = 8'hC9;
    buff [16'h01_02] = 8'hFB;
    buff [16'h01_03] = 8'hE4;
    buff [16'h01_04] = 8'hCA;
    buff [16'h01_05] = 8'hFC;
    buff [16'h01_06] = 8'hE8;
    buff [16'h01_07] = 8'h30;
    buff [16'h01_08] = 8'hE3;
    buff [16'h01_09] = 8'h05;
    buff [16'h01_0a] = 8'hE4;
    buff [16'h01_0b] = 8'hC9;
    buff [16'h01_0c] = 8'hCA;
    buff [16'h01_0d] = 8'hCB;
    buff [16'h01_0e] = 8'hFC;
    buff [16'h01_0f] = 8'hE8;
    buff [16'h01_10] = 8'h54;
    buff [16'h01_11] = 8'h07;
    buff [16'h01_12] = 8'h60;
    buff [16'h01_13] = 8'h10;
    buff [16'h01_14] = 8'hF8;
    buff [16'h01_15] = 8'hC3;
    buff [16'h01_16] = 8'hE9;
    buff [16'h01_17] = 8'h13;
    buff [16'h01_18] = 8'hF9;
    buff [16'h01_19] = 8'hEA;
    buff [16'h01_1a] = 8'h13;
    buff [16'h01_1b] = 8'hFA;
    buff [16'h01_1c] = 8'hEB;
    buff [16'h01_1d] = 8'h13;
    buff [16'h01_1e] = 8'hFB;
    buff [16'h01_1f] = 8'hEC;
    buff [16'h01_20] = 8'h13;
    buff [16'h01_21] = 8'hFC;
    buff [16'h01_22] = 8'hD8;
    buff [16'h01_23] = 8'hF1;
    buff [16'h01_24] = 8'h30;
    buff [16'h01_25] = 8'hF5;
    buff [16'h01_26] = 8'h2F;
    buff [16'h01_27] = 8'hC3;
    buff [16'h01_28] = 8'hE4;
    buff [16'h01_29] = 8'h9C;
    buff [16'h01_2a] = 8'hFC;
    buff [16'h01_2b] = 8'hEF;
    buff [16'h01_2c] = 8'h9B;
    buff [16'h01_2d] = 8'hFF;
    buff [16'h01_2e] = 8'hEE;
    buff [16'h01_2f] = 8'h9A;
    buff [16'h01_30] = 8'hFE;
    buff [16'h01_31] = 8'hED;
    buff [16'h01_32] = 8'h99;
    buff [16'h01_33] = 8'hFD;
    buff [16'h01_34] = 8'hD0;
    buff [16'h01_35] = 8'hE0;
    buff [16'h01_36] = 8'hFB;
    buff [16'h01_37] = 8'hEF;
    buff [16'h01_38] = 8'h4E;
    buff [16'h01_39] = 8'h4D;
    buff [16'h01_3a] = 8'h4C;
    buff [16'h01_3b] = 8'h70;
    buff [16'h01_3c] = 8'h12;
    buff [16'h01_3d] = 8'h22;
    buff [16'h01_3e] = 8'hDB;
    buff [16'h01_3f] = 8'h03;
    buff [16'h01_40] = 8'h02;
    buff [16'h01_41] = 8'h02;
    buff [16'h01_42] = 8'hF3;
    buff [16'h01_43] = 8'hEC;
    buff [16'h01_44] = 8'h2C;
    buff [16'h01_45] = 8'hFC;
    buff [16'h01_46] = 8'hEF;
    buff [16'h01_47] = 8'h33;
    buff [16'h01_48] = 8'hFF;
    buff [16'h01_49] = 8'hEE;
    buff [16'h01_4a] = 8'h33;
    buff [16'h01_4b] = 8'hFE;
    buff [16'h01_4c] = 8'hED;
    buff [16'h01_4d] = 8'h33;
    buff [16'h01_4e] = 8'hFD;
    buff [16'h01_4f] = 8'hED;
    buff [16'h01_50] = 8'h30;
    buff [16'h01_51] = 8'hE7;
    buff [16'h01_52] = 8'hEB;
    buff [16'h01_53] = 8'h02;
    buff [16'h01_54] = 8'h02;
    buff [16'h01_55] = 8'hCE;
    buff [16'h01_56] = 8'hEF;
    buff [16'h01_57] = 8'h2B;
    buff [16'h01_58] = 8'hFF;
    buff [16'h01_59] = 8'hEE;
    buff [16'h01_5a] = 8'h3A;
    buff [16'h01_5b] = 8'hFE;
    buff [16'h01_5c] = 8'hED;
    buff [16'h01_5d] = 8'h39;
    buff [16'h01_5e] = 8'hFD;
    buff [16'h01_5f] = 8'hD0;
    buff [16'h01_60] = 8'hE0;
    buff [16'h01_61] = 8'hFB;
    buff [16'h01_62] = 8'h50;
    buff [16'h01_63] = 8'h13;
    buff [16'h01_64] = 8'h0B;
    buff [16'h01_65] = 8'hBB;
    buff [16'h01_66] = 8'h00;
    buff [16'h01_67] = 8'h03;
    buff [16'h01_68] = 8'h02;
    buff [16'h01_69] = 8'h02;
    buff [16'h01_6a] = 8'hF6;
    buff [16'h01_6b] = 8'hED;
    buff [16'h01_6c] = 8'h13;
    buff [16'h01_6d] = 8'hFD;
    buff [16'h01_6e] = 8'hEE;
    buff [16'h01_6f] = 8'h13;
    buff [16'h01_70] = 8'hFE;
    buff [16'h01_71] = 8'hEF;
    buff [16'h01_72] = 8'h13;
    buff [16'h01_73] = 8'hFF;
    buff [16'h01_74] = 8'hEC;
    buff [16'h01_75] = 8'h13;
    buff [16'h01_76] = 8'hFC;
    buff [16'h01_77] = 8'h02;
    buff [16'h01_78] = 8'h02;
    buff [16'h01_79] = 8'hCE;
    buff [16'h01_7a] = 8'hEC;
    buff [16'h01_7b] = 8'h4D;
    buff [16'h01_7c] = 8'h60;
    buff [16'h01_7d] = 8'h11;
    buff [16'h01_7e] = 8'hE8;
    buff [16'h01_7f] = 8'h49;
    buff [16'h01_80] = 8'h70;
    buff [16'h01_81] = 8'h17;
    buff [16'h01_82] = 8'hED;
    buff [16'h01_83] = 8'h33;
    buff [16'h01_84] = 8'hEC;
    buff [16'h01_85] = 8'h33;
    buff [16'h01_86] = 8'h04;
    buff [16'h01_87] = 8'h60;
    buff [16'h01_88] = 8'h0D;
    buff [16'h01_89] = 8'hE4;
    buff [16'h01_8a] = 8'hFC;
    buff [16'h01_8b] = 8'hFF;
    buff [16'h01_8c] = 8'hFE;
    buff [16'h01_8d] = 8'hFD;
    buff [16'h01_8e] = 8'h22;
    buff [16'h01_8f] = 8'hE9;
    buff [16'h01_90] = 8'h33;
    buff [16'h01_91] = 8'hE8;
    buff [16'h01_92] = 8'h33;
    buff [16'h01_93] = 8'h04;
    buff [16'h01_94] = 8'h70;
    buff [16'h01_95] = 8'hF8;
    buff [16'h01_96] = 8'h02;
    buff [16'h01_97] = 8'h02;
    buff [16'h01_98] = 8'hEC;
    buff [16'h01_99] = 8'h12;
    buff [16'h01_9a] = 8'h02;
    buff [16'h01_9b] = 8'hB7;
    buff [16'h01_9c] = 8'h58;
    buff [16'h01_9d] = 8'h04;
    buff [16'h01_9e] = 8'h60;
    buff [16'h01_9f] = 8'h09;
    buff [16'h01_a0] = 8'hE4;
    buff [16'h01_a1] = 8'hCC;
    buff [16'h01_a2] = 8'h24;
    buff [16'h01_a3] = 8'h81;
    buff [16'h01_a4] = 8'h50;
    buff [16'h01_a5] = 8'h06;
    buff [16'h01_a6] = 8'h28;
    buff [16'h01_a7] = 8'h50;
    buff [16'h01_a8] = 8'h09;
    buff [16'h01_a9] = 8'h02;
    buff [16'h01_aa] = 8'h02;
    buff [16'h01_ab] = 8'hF6;
    buff [16'h01_ac] = 8'h28;
    buff [16'h01_ad] = 8'h40;
    buff [16'h01_ae] = 8'h03;
    buff [16'h01_af] = 8'h02;
    buff [16'h01_b0] = 8'h02;
    buff [16'h01_b1] = 8'hF3;
    buff [16'h01_b2] = 8'hC0;
    buff [16'h01_b3] = 8'hE0;
    buff [16'h01_b4] = 8'hEB;
    buff [16'h01_b5] = 8'h4A;
    buff [16'h01_b6] = 8'h70;
    buff [16'h01_b7] = 8'h44;
    buff [16'h01_b8] = 8'hB9;
    buff [16'h01_b9] = 8'h80;
    buff [16'h01_ba] = 8'h06;
    buff [16'h01_bb] = 8'hD0;
    buff [16'h01_bc] = 8'hE0;
    buff [16'h01_bd] = 8'hFB;
    buff [16'h01_be] = 8'h02;
    buff [16'h01_bf] = 8'h02;
    buff [16'h01_c0] = 8'hE2;
    buff [16'h01_c1] = 8'hEF;
    buff [16'h01_c2] = 8'h4E;
    buff [16'h01_c3] = 8'h70;
    buff [16'h01_c4] = 8'h1C;
    buff [16'h01_c5] = 8'hBD;
    buff [16'h01_c6] = 8'h80;
    buff [16'h01_c7] = 8'h08;
    buff [16'h01_c8] = 8'hEB;
    buff [16'h01_c9] = 8'hFF;
    buff [16'h01_ca] = 8'hEA;
    buff [16'h01_cb] = 8'hFE;
    buff [16'h01_cc] = 8'hE9;
    buff [16'h01_cd] = 8'hFD;
    buff [16'h01_ce] = 8'h80;
    buff [16'h01_cf] = 8'hEB;
    buff [16'h01_d0] = 8'hE9;
    buff [16'h01_d1] = 8'h8D;
    buff [16'h01_d2] = 8'hF0;
    buff [16'h01_d3] = 8'hA4;
    buff [16'h01_d4] = 8'hFE;
    buff [16'h01_d5] = 8'hE5;
    buff [16'h01_d6] = 8'hF0;
    buff [16'h01_d7] = 8'h02;
    buff [16'h01_d8] = 8'h02;
    buff [16'h01_d9] = 8'h63;
    buff [16'h01_da] = 8'hE9;
    buff [16'h01_db] = 8'hCD;
    buff [16'h01_dc] = 8'hF9;
    buff [16'h01_dd] = 8'hEA;
    buff [16'h01_de] = 8'hFE;
    buff [16'h01_df] = 8'hEB;
    buff [16'h01_e0] = 8'hFF;
    buff [16'h01_e1] = 8'hEF;
    buff [16'h01_e2] = 8'h89;
    buff [16'h01_e3] = 8'hF0;
    buff [16'h01_e4] = 8'hA4;
    buff [16'h01_e5] = 8'hFC;
    buff [16'h01_e6] = 8'hE5;
    buff [16'h01_e7] = 8'hF0;
    buff [16'h01_e8] = 8'hCE;
    buff [16'h01_e9] = 8'h89;
    buff [16'h01_ea] = 8'hF0;
    buff [16'h01_eb] = 8'hA4;
    buff [16'h01_ec] = 8'h2E;
    buff [16'h01_ed] = 8'hFF;
    buff [16'h01_ee] = 8'hE4;
    buff [16'h01_ef] = 8'h35;
    buff [16'h01_f0] = 8'hF0;
    buff [16'h01_f1] = 8'hCD;
    buff [16'h01_f2] = 8'h89;
    buff [16'h01_f3] = 8'hF0;
    buff [16'h01_f4] = 8'hA4;
    buff [16'h01_f5] = 8'h2D;
    buff [16'h01_f6] = 8'hFE;
    buff [16'h01_f7] = 8'hE4;
    buff [16'h01_f8] = 8'h35;
    buff [16'h01_f9] = 8'hF0;
    buff [16'h01_fa] = 8'h80;
    buff [16'h01_fb] = 8'h67;
    buff [16'h01_fc] = 8'hEF;
    buff [16'h01_fd] = 8'h4E;
    buff [16'h01_fe] = 8'h70;
    buff [16'h01_ff] = 8'h05;
    buff [16'h02_00] = 8'hBD;
    buff [16'h02_01] = 8'h80;
    buff [16'h02_02] = 8'hD7;
    buff [16'h02_03] = 8'h80;
    buff [16'h02_04] = 8'hC3;
    buff [16'h02_05] = 8'hEF;
    buff [16'h02_06] = 8'h8B;
    buff [16'h02_07] = 8'hF0;
    buff [16'h02_08] = 8'hA4;
    buff [16'h02_09] = 8'hAC;
    buff [16'h02_0a] = 8'hF0;
    buff [16'h02_0b] = 8'hEE;
    buff [16'h02_0c] = 8'h8B;
    buff [16'h02_0d] = 8'hF0;
    buff [16'h02_0e] = 8'hA4;
    buff [16'h02_0f] = 8'h2C;
    buff [16'h02_10] = 8'hFC;
    buff [16'h02_11] = 8'hE4;
    buff [16'h02_12] = 8'h35;
    buff [16'h02_13] = 8'hF0;
    buff [16'h02_14] = 8'hF8;
    buff [16'h02_15] = 8'hEF;
    buff [16'h02_16] = 8'h8A;
    buff [16'h02_17] = 8'hF0;
    buff [16'h02_18] = 8'hA4;
    buff [16'h02_19] = 8'h2C;
    buff [16'h02_1a] = 8'hE5;
    buff [16'h02_1b] = 8'hF0;
    buff [16'h02_1c] = 8'h38;
    buff [16'h02_1d] = 8'hFC;
    buff [16'h02_1e] = 8'hE4;
    buff [16'h02_1f] = 8'h33;
    buff [16'h02_20] = 8'hCB;
    buff [16'h02_21] = 8'h8D;
    buff [16'h02_22] = 8'hF0;
    buff [16'h02_23] = 8'hA4;
    buff [16'h02_24] = 8'h2C;
    buff [16'h02_25] = 8'hFC;
    buff [16'h02_26] = 8'hE5;
    buff [16'h02_27] = 8'hF0;
    buff [16'h02_28] = 8'h3B;
    buff [16'h02_29] = 8'hF8;
    buff [16'h02_2a] = 8'hEE;
    buff [16'h02_2b] = 8'h8A;
    buff [16'h02_2c] = 8'hF0;
    buff [16'h02_2d] = 8'hA4;
    buff [16'h02_2e] = 8'h2C;
    buff [16'h02_2f] = 8'hFC;
    buff [16'h02_30] = 8'hE5;
    buff [16'h02_31] = 8'hF0;
    buff [16'h02_32] = 8'h38;
    buff [16'h02_33] = 8'hF8;
    buff [16'h02_34] = 8'hE4;
    buff [16'h02_35] = 8'h33;
    buff [16'h02_36] = 8'hCF;
    buff [16'h02_37] = 8'h89;
    buff [16'h02_38] = 8'hF0;
    buff [16'h02_39] = 8'hA4;
    buff [16'h02_3a] = 8'h2C;
    buff [16'h02_3b] = 8'hFC;
    buff [16'h02_3c] = 8'hE5;
    buff [16'h02_3d] = 8'hF0;
    buff [16'h02_3e] = 8'h38;
    buff [16'h02_3f] = 8'hCF;
    buff [16'h02_40] = 8'h34;
    buff [16'h02_41] = 8'h00;
    buff [16'h02_42] = 8'hCE;
    buff [16'h02_43] = 8'h89;
    buff [16'h02_44] = 8'hF0;
    buff [16'h02_45] = 8'hA4;
    buff [16'h02_46] = 8'h2F;
    buff [16'h02_47] = 8'hFF;
    buff [16'h02_48] = 8'hE5;
    buff [16'h02_49] = 8'hF0;
    buff [16'h02_4a] = 8'h3E;
    buff [16'h02_4b] = 8'hFE;
    buff [16'h02_4c] = 8'hE4;
    buff [16'h02_4d] = 8'h33;
    buff [16'h02_4e] = 8'hC9;
    buff [16'h02_4f] = 8'h8D;
    buff [16'h02_50] = 8'hF0;
    buff [16'h02_51] = 8'hA4;
    buff [16'h02_52] = 8'h2E;
    buff [16'h02_53] = 8'hFE;
    buff [16'h02_54] = 8'hE5;
    buff [16'h02_55] = 8'hF0;
    buff [16'h02_56] = 8'h39;
    buff [16'h02_57] = 8'hCD;
    buff [16'h02_58] = 8'h8A;
    buff [16'h02_59] = 8'hF0;
    buff [16'h02_5a] = 8'hA4;
    buff [16'h02_5b] = 8'h2F;
    buff [16'h02_5c] = 8'hFF;
    buff [16'h02_5d] = 8'hE5;
    buff [16'h02_5e] = 8'hF0;
    buff [16'h02_5f] = 8'h3E;
    buff [16'h02_60] = 8'hFE;
    buff [16'h02_61] = 8'hE4;
    buff [16'h02_62] = 8'h3D;
    buff [16'h02_63] = 8'hFD;
    buff [16'h02_64] = 8'h33;
    buff [16'h02_65] = 8'hD0;
    buff [16'h02_66] = 8'hE0;
    buff [16'h02_67] = 8'hFB;
    buff [16'h02_68] = 8'h50;
    buff [16'h02_69] = 8'h07;
    buff [16'h02_6a] = 8'h0B;
    buff [16'h02_6b] = 8'hBB;
    buff [16'h02_6c] = 8'h00;
    buff [16'h02_6d] = 8'h0F;
    buff [16'h02_6e] = 8'h02;
    buff [16'h02_6f] = 8'h02;
    buff [16'h02_70] = 8'hF6;
    buff [16'h02_71] = 8'hEC;
    buff [16'h02_72] = 8'h2C;
    buff [16'h02_73] = 8'hFC;
    buff [16'h02_74] = 8'hEF;
    buff [16'h02_75] = 8'h33;
    buff [16'h02_76] = 8'hFF;
    buff [16'h02_77] = 8'hEE;
    buff [16'h02_78] = 8'h33;
    buff [16'h02_79] = 8'hFE;
    buff [16'h02_7a] = 8'hED;
    buff [16'h02_7b] = 8'h33;
    buff [16'h02_7c] = 8'hFD;
    buff [16'h02_7d] = 8'h02;
    buff [16'h02_7e] = 8'h02;
    buff [16'h02_7f] = 8'hCE;
    buff [16'h02_80] = 8'hED;
    buff [16'h02_81] = 8'hD2;
    buff [16'h02_82] = 8'hE7;
    buff [16'h02_83] = 8'hCD;
    buff [16'h02_84] = 8'h33;
    buff [16'h02_85] = 8'hEC;
    buff [16'h02_86] = 8'h33;
    buff [16'h02_87] = 8'h92;
    buff [16'h02_88] = 8'hD5;
    buff [16'h02_89] = 8'h24;
    buff [16'h02_8a] = 8'h81;
    buff [16'h02_8b] = 8'h40;
    buff [16'h02_8c] = 8'h06;
    buff [16'h02_8d] = 8'hE4;
    buff [16'h02_8e] = 8'hFF;
    buff [16'h02_8f] = 8'hFE;
    buff [16'h02_90] = 8'hFD;
    buff [16'h02_91] = 8'hFC;
    buff [16'h02_92] = 8'h22;
    buff [16'h02_93] = 8'hFC;
    buff [16'h02_94] = 8'hE4;
    buff [16'h02_95] = 8'hCF;
    buff [16'h02_96] = 8'hCE;
    buff [16'h02_97] = 8'hCD;
    buff [16'h02_98] = 8'hCC;
    buff [16'h02_99] = 8'h24;
    buff [16'h02_9a] = 8'hE0;
    buff [16'h02_9b] = 8'h50;
    buff [16'h02_9c] = 8'h11;
    buff [16'h02_9d] = 8'h74;
    buff [16'h02_9e] = 8'hFF;
    buff [16'h02_9f] = 8'h80;
    buff [16'h02_a0] = 8'hED;
    buff [16'h02_a1] = 8'hC3;
    buff [16'h02_a2] = 8'hCC;
    buff [16'h02_a3] = 8'h13;
    buff [16'h02_a4] = 8'hCC;
    buff [16'h02_a5] = 8'hCD;
    buff [16'h02_a6] = 8'h13;
    buff [16'h02_a7] = 8'hCD;
    buff [16'h02_a8] = 8'hCE;
    buff [16'h02_a9] = 8'h13;
    buff [16'h02_aa] = 8'hCE;
    buff [16'h02_ab] = 8'hCF;
    buff [16'h02_ac] = 8'h13;
    buff [16'h02_ad] = 8'hCF;
    buff [16'h02_ae] = 8'h04;
    buff [16'h02_af] = 8'h70;
    buff [16'h02_b0] = 8'hF0;
    buff [16'h02_b1] = 8'h30;
    buff [16'h02_b2] = 8'hD5;
    buff [16'h02_b3] = 8'hDE;
    buff [16'h02_b4] = 8'h02;
    buff [16'h02_b5] = 8'h03;
    buff [16'h02_b6] = 8'h9C;
    buff [16'h02_b7] = 8'hE9;
    buff [16'h02_b8] = 8'hD2;
    buff [16'h02_b9] = 8'hE7;
    buff [16'h02_ba] = 8'hC9;
    buff [16'h02_bb] = 8'h33;
    buff [16'h02_bc] = 8'hE8;
    buff [16'h02_bd] = 8'h33;
    buff [16'h02_be] = 8'hF8;
    buff [16'h02_bf] = 8'h92;
    buff [16'h02_c0] = 8'hD5;
    buff [16'h02_c1] = 8'hED;
    buff [16'h02_c2] = 8'hD2;
    buff [16'h02_c3] = 8'hE7;
    buff [16'h02_c4] = 8'hCD;
    buff [16'h02_c5] = 8'h33;
    buff [16'h02_c6] = 8'hEC;
    buff [16'h02_c7] = 8'h33;
    buff [16'h02_c8] = 8'hFC;
    buff [16'h02_c9] = 8'h50;
    buff [16'h02_ca] = 8'h02;
    buff [16'h02_cb] = 8'hB2;
    buff [16'h02_cc] = 8'hD5;
    buff [16'h02_cd] = 8'h22;
    buff [16'h02_ce] = 8'hEC;
    buff [16'h02_cf] = 8'h30;
    buff [16'h02_d0] = 8'hE7;
    buff [16'h02_d1] = 8'h10;
    buff [16'h02_d2] = 8'h0F;
    buff [16'h02_d3] = 8'hBF;
    buff [16'h02_d4] = 8'h00;
    buff [16'h02_d5] = 8'h0C;
    buff [16'h02_d6] = 8'h0E;
    buff [16'h02_d7] = 8'hBE;
    buff [16'h02_d8] = 8'h00;
    buff [16'h02_d9] = 8'h08;
    buff [16'h02_da] = 8'h0D;
    buff [16'h02_db] = 8'hBD;
    buff [16'h02_dc] = 8'h00;
    buff [16'h02_dd] = 8'h04;
    buff [16'h02_de] = 8'h0B;
    buff [16'h02_df] = 8'hEB;
    buff [16'h02_e0] = 8'h60;
    buff [16'h02_e1] = 8'h14;
    buff [16'h02_e2] = 8'hA2;
    buff [16'h02_e3] = 8'hD5;
    buff [16'h02_e4] = 8'hEB;
    buff [16'h02_e5] = 8'h13;
    buff [16'h02_e6] = 8'hFC;
    buff [16'h02_e7] = 8'hED;
    buff [16'h02_e8] = 8'h92;
    buff [16'h02_e9] = 8'hE7;
    buff [16'h02_ea] = 8'hFD;
    buff [16'h02_eb] = 8'h22;
    buff [16'h02_ec] = 8'h74;
    buff [16'h02_ed] = 8'hFF;
    buff [16'h02_ee] = 8'hFC;
    buff [16'h02_ef] = 8'hFD;
    buff [16'h02_f0] = 8'hFE;
    buff [16'h02_f1] = 8'hFF;
    buff [16'h02_f2] = 8'h22;
    buff [16'h02_f3] = 8'hE4;
    buff [16'h02_f4] = 8'h80;
    buff [16'h02_f5] = 8'hF8;
    buff [16'h02_f6] = 8'hA2;
    buff [16'h02_f7] = 8'hD5;
    buff [16'h02_f8] = 8'h74;
    buff [16'h02_f9] = 8'hFF;
    buff [16'h02_fa] = 8'h13;
    buff [16'h02_fb] = 8'hFC;
    buff [16'h02_fc] = 8'h7D;
    buff [16'h02_fd] = 8'h80;
    buff [16'h02_fe] = 8'h80;
    buff [16'h02_ff] = 8'hF0;
    buff [16'h03_00] = 8'h02;
    buff [16'h03_01] = 8'h02;
    buff [16'h03_02] = 8'hF6;
    buff [16'h03_03] = 8'hEC;
    buff [16'h03_04] = 8'h5D;
    buff [16'h03_05] = 8'h04;
    buff [16'h03_06] = 8'h60;
    buff [16'h03_07] = 8'h05;
    buff [16'h03_08] = 8'hE8;
    buff [16'h03_09] = 8'h59;
    buff [16'h03_0a] = 8'h04;
    buff [16'h03_0b] = 8'h70;
    buff [16'h03_0c] = 8'h03;
    buff [16'h03_0d] = 8'h02;
    buff [16'h03_0e] = 8'h02;
    buff [16'h03_0f] = 8'hEC;
    buff [16'h03_10] = 8'h12;
    buff [16'h03_11] = 8'h02;
    buff [16'h03_12] = 8'hB7;
    buff [16'h03_13] = 8'h58;
    buff [16'h03_14] = 8'h04;
    buff [16'h03_15] = 8'h60;
    buff [16'h03_16] = 8'hF6;
    buff [16'h03_17] = 8'hEC;
    buff [16'h03_18] = 8'h48;
    buff [16'h03_19] = 8'h60;
    buff [16'h03_1a] = 8'hF2;
    buff [16'h03_1b] = 8'hEC;
    buff [16'h03_1c] = 8'h70;
    buff [16'h03_1d] = 8'h04;
    buff [16'h03_1e] = 8'hFD;
    buff [16'h03_1f] = 8'hFE;
    buff [16'h03_20] = 8'hFF;
    buff [16'h03_21] = 8'h22;
    buff [16'h03_22] = 8'hC8;
    buff [16'h03_23] = 8'h24;
    buff [16'h03_24] = 8'h81;
    buff [16'h03_25] = 8'hC8;
    buff [16'h03_26] = 8'h50;
    buff [16'h03_27] = 8'h07;
    buff [16'h03_28] = 8'hC3;
    buff [16'h03_29] = 8'h98;
    buff [16'h03_2a] = 8'h50;
    buff [16'h03_2b] = 8'h06;
    buff [16'h03_2c] = 8'h02;
    buff [16'h03_2d] = 8'h02;
    buff [16'h03_2e] = 8'hF3;
    buff [16'h03_2f] = 8'h98;
    buff [16'h03_30] = 8'h50;
    buff [16'h03_31] = 8'hCE;
    buff [16'h03_32] = 8'hF5;
    buff [16'h03_33] = 8'h82;
    buff [16'h03_34] = 8'hE9;
    buff [16'h03_35] = 8'h29;
    buff [16'h03_36] = 8'h4B;
    buff [16'h03_37] = 8'h4A;
    buff [16'h03_38] = 8'h70;
    buff [16'h03_39] = 8'h05;
    buff [16'h03_3a] = 8'hAB;
    buff [16'h03_3b] = 8'h82;
    buff [16'h03_3c] = 8'h02;
    buff [16'h03_3d] = 8'h02;
    buff [16'h03_3e] = 8'hE2;
    buff [16'h03_3f] = 8'h75;
    buff [16'h03_40] = 8'hF0;
    buff [16'h03_41] = 8'h00;
    buff [16'h03_42] = 8'h7C;
    buff [16'h03_43] = 8'h1A;
    buff [16'h03_44] = 8'h78;
    buff [16'h03_45] = 8'h80;
    buff [16'h03_46] = 8'hC3;
    buff [16'h03_47] = 8'hEF;
    buff [16'h03_48] = 8'h9B;
    buff [16'h03_49] = 8'hEE;
    buff [16'h03_4a] = 8'h9A;
    buff [16'h03_4b] = 8'hED;
    buff [16'h03_4c] = 8'h99;
    buff [16'h03_4d] = 8'h40;
    buff [16'h03_4e] = 8'h0D;
    buff [16'h03_4f] = 8'hC3;
    buff [16'h03_50] = 8'hEF;
    buff [16'h03_51] = 8'h9B;
    buff [16'h03_52] = 8'hFF;
    buff [16'h03_53] = 8'hEE;
    buff [16'h03_54] = 8'h9A;
    buff [16'h03_55] = 8'hFE;
    buff [16'h03_56] = 8'hED;
    buff [16'h03_57] = 8'h99;
    buff [16'h03_58] = 8'hFD;
    buff [16'h03_59] = 8'hE8;
    buff [16'h03_5a] = 8'h42;
    buff [16'h03_5b] = 8'hF0;
    buff [16'h03_5c] = 8'hDC;
    buff [16'h03_5d] = 8'h23;
    buff [16'h03_5e] = 8'hAC;
    buff [16'h03_5f] = 8'hF0;
    buff [16'h03_60] = 8'hD0;
    buff [16'h03_61] = 8'hE0;
    buff [16'h03_62] = 8'hFF;
    buff [16'h03_63] = 8'hD0;
    buff [16'h03_64] = 8'hE0;
    buff [16'h03_65] = 8'hFE;
    buff [16'h03_66] = 8'hD0;
    buff [16'h03_67] = 8'hE0;
    buff [16'h03_68] = 8'hFD;
    buff [16'h03_69] = 8'hAB;
    buff [16'h03_6a] = 8'h82;
    buff [16'h03_6b] = 8'h20;
    buff [16'h03_6c] = 8'hE7;
    buff [16'h03_6d] = 8'h10;
    buff [16'h03_6e] = 8'h1B;
    buff [16'h03_6f] = 8'hEB;
    buff [16'h03_70] = 8'h60;
    buff [16'h03_71] = 8'hBA;
    buff [16'h03_72] = 8'hEC;
    buff [16'h03_73] = 8'h2C;
    buff [16'h03_74] = 8'hFC;
    buff [16'h03_75] = 8'hEF;
    buff [16'h03_76] = 8'h33;
    buff [16'h03_77] = 8'hFF;
    buff [16'h03_78] = 8'hEE;
    buff [16'h03_79] = 8'h33;
    buff [16'h03_7a] = 8'hFE;
    buff [16'h03_7b] = 8'hED;
    buff [16'h03_7c] = 8'h33;
    buff [16'h03_7d] = 8'hFD;
    buff [16'h03_7e] = 8'h02;
    buff [16'h03_7f] = 8'h02;
    buff [16'h03_80] = 8'hCE;
    buff [16'h03_81] = 8'hE8;
    buff [16'h03_82] = 8'h03;
    buff [16'h03_83] = 8'hF8;
    buff [16'h03_84] = 8'h30;
    buff [16'h03_85] = 8'hE7;
    buff [16'h03_86] = 8'h05;
    buff [16'h03_87] = 8'hC0;
    buff [16'h03_88] = 8'hF0;
    buff [16'h03_89] = 8'h75;
    buff [16'h03_8a] = 8'hF0;
    buff [16'h03_8b] = 8'h00;
    buff [16'h03_8c] = 8'hEF;
    buff [16'h03_8d] = 8'h2F;
    buff [16'h03_8e] = 8'hFF;
    buff [16'h03_8f] = 8'hEE;
    buff [16'h03_90] = 8'h33;
    buff [16'h03_91] = 8'hFE;
    buff [16'h03_92] = 8'hED;
    buff [16'h03_93] = 8'h33;
    buff [16'h03_94] = 8'hFD;
    buff [16'h03_95] = 8'h40;
    buff [16'h03_96] = 8'hB8;
    buff [16'h03_97] = 8'h30;
    buff [16'h03_98] = 8'hE7;
    buff [16'h03_99] = 8'hC2;
    buff [16'h03_9a] = 8'h80;
    buff [16'h03_9b] = 8'hAA;
    buff [16'h03_9c] = 8'hC3;
    buff [16'h03_9d] = 8'hE4;
    buff [16'h03_9e] = 8'h9F;
    buff [16'h03_9f] = 8'hFF;
    buff [16'h03_a0] = 8'hE4;
    buff [16'h03_a1] = 8'h9E;
    buff [16'h03_a2] = 8'hFE;
    buff [16'h03_a3] = 8'hE4;
    buff [16'h03_a4] = 8'h9D;
    buff [16'h03_a5] = 8'hFD;
    buff [16'h03_a6] = 8'hE4;
    buff [16'h03_a7] = 8'h9C;
    buff [16'h03_a8] = 8'hFC;
    buff [16'h03_a9] = 8'h22;
    buff [16'h03_aa] = 8'h02;
    buff [16'h03_ab] = 8'h02;
    buff [16'h03_ac] = 8'hEC;
    buff [16'h03_ad] = 8'h22;
    buff [16'h03_ae] = 8'hED;
    buff [16'h03_af] = 8'hA2;
    buff [16'h03_b0] = 8'hE7;
    buff [16'h03_b1] = 8'hD2;
    buff [16'h03_b2] = 8'hE7;
    buff [16'h03_b3] = 8'hF9;
    buff [16'h03_b4] = 8'hEC;
    buff [16'h03_b5] = 8'h33;
    buff [16'h03_b6] = 8'h40;
    buff [16'h03_b7] = 8'hF2;
    buff [16'h03_b8] = 8'h60;
    buff [16'h03_b9] = 8'hF3;
    buff [16'h03_ba] = 8'hB4;
    buff [16'h03_bb] = 8'hFF;
    buff [16'h03_bc] = 8'h08;
    buff [16'h03_bd] = 8'hED;
    buff [16'h03_be] = 8'h54;
    buff [16'h03_bf] = 8'h7F;
    buff [16'h03_c0] = 8'h70;
    buff [16'h03_c1] = 8'hE8;
    buff [16'h03_c2] = 8'h02;
    buff [16'h03_c3] = 8'h02;
    buff [16'h03_c4] = 8'hF6;
    buff [16'h03_c5] = 8'hF8;
    buff [16'h03_c6] = 8'h24;
    buff [16'h03_c7] = 8'h81;
    buff [16'h03_c8] = 8'hC2;
    buff [16'h03_c9] = 8'hE0;
    buff [16'h03_ca] = 8'hC0;
    buff [16'h03_cb] = 8'hE0;
    buff [16'h03_cc] = 8'hF4;
    buff [16'h03_cd] = 8'h04;
    buff [16'h03_ce] = 8'h28;
    buff [16'h03_cf] = 8'hFA;
    buff [16'h03_d0] = 8'hC3;
    buff [16'h03_d1] = 8'h13;
    buff [16'h03_d2] = 8'hFC;
    buff [16'h03_d3] = 8'hED;
    buff [16'h03_d4] = 8'h92;
    buff [16'h03_d5] = 8'hE7;
    buff [16'h03_d6] = 8'hFD;
    buff [16'h03_d7] = 8'h8C;
    buff [16'h03_d8] = 8'h18;
    buff [16'h03_d9] = 8'h8D;
    buff [16'h03_da] = 8'h19;
    buff [16'h03_db] = 8'h8E;
    buff [16'h03_dc] = 8'h1A;
    buff [16'h03_dd] = 8'h8F;
    buff [16'h03_de] = 8'h1B;
    buff [16'h03_df] = 8'hEE;
    buff [16'h03_e0] = 8'hA2;
    buff [16'h03_e1] = 8'hE7;
    buff [16'h03_e2] = 8'hE9;
    buff [16'h03_e3] = 8'hBA;
    buff [16'h03_e4] = 8'h7F;
    buff [16'h03_e5] = 8'h02;
    buff [16'h03_e6] = 8'hC3;
    buff [16'h03_e7] = 8'h13;
    buff [16'h03_e8] = 8'h34;
    buff [16'h03_e9] = 8'h00;
    buff [16'h03_ea] = 8'h94;
    buff [16'h03_eb] = 8'h00;
    buff [16'h03_ec] = 8'hFA;
    buff [16'h03_ed] = 8'h75;
    buff [16'h03_ee] = 8'hF0;
    buff [16'h03_ef] = 8'h91;
    buff [16'h03_f0] = 8'hA4;
    buff [16'h03_f1] = 8'hE5;
    buff [16'h03_f2] = 8'hF0;
    buff [16'h03_f3] = 8'h13;
    buff [16'h03_f4] = 8'hF4;
    buff [16'h03_f5] = 8'h94;
    buff [16'h03_f6] = 8'hFE;
    buff [16'h03_f7] = 8'h8A;
    buff [16'h03_f8] = 8'hF0;
    buff [16'h03_f9] = 8'hA4;
    buff [16'h03_fa] = 8'h33;
    buff [16'h03_fb] = 8'hE5;
    buff [16'h03_fc] = 8'hF0;
    buff [16'h03_fd] = 8'h33;
    buff [16'h03_fe] = 8'h24;
    buff [16'h03_ff] = 8'h8C;
    buff [16'h04_00] = 8'hD3;
    buff [16'h04_01] = 8'h13;
    buff [16'h04_02] = 8'hFD;
    buff [16'h04_03] = 8'hE4;
    buff [16'h04_04] = 8'h92;
    buff [16'h04_05] = 8'hE7;
    buff [16'h04_06] = 8'hFE;
    buff [16'h04_07] = 8'h7F;
    buff [16'h04_08] = 8'h00;
    buff [16'h04_09] = 8'h7C;
    buff [16'h04_0a] = 8'h3F;
    buff [16'h04_0b] = 8'h75;
    buff [16'h04_0c] = 8'h83;
    buff [16'h04_0d] = 8'h02;
    buff [16'h04_0e] = 8'hEC;
    buff [16'h04_0f] = 8'hC0;
    buff [16'h04_10] = 8'hE0;
    buff [16'h04_11] = 8'hF8;
    buff [16'h04_12] = 8'hED;
    buff [16'h04_13] = 8'hC0;
    buff [16'h04_14] = 8'hE0;
    buff [16'h04_15] = 8'hF9;
    buff [16'h04_16] = 8'hEE;
    buff [16'h04_17] = 8'hC0;
    buff [16'h04_18] = 8'hE0;
    buff [16'h04_19] = 8'hFA;
    buff [16'h04_1a] = 8'hEF;
    buff [16'h04_1b] = 8'hC0;
    buff [16'h04_1c] = 8'hE0;
    buff [16'h04_1d] = 8'hFB;
    buff [16'h04_1e] = 8'hAC;
    buff [16'h04_1f] = 8'h18;
    buff [16'h04_20] = 8'hAD;
    buff [16'h04_21] = 8'h19;
    buff [16'h04_22] = 8'hAE;
    buff [16'h04_23] = 8'h1A;
    buff [16'h04_24] = 8'hAF;
    buff [16'h04_25] = 8'h1B;
    buff [16'h04_26] = 8'h12;
    buff [16'h04_27] = 8'h03;
    buff [16'h04_28] = 8'h03;
    buff [16'h04_29] = 8'hD0;
    buff [16'h04_2a] = 8'hE0;
    buff [16'h04_2b] = 8'hFB;
    buff [16'h04_2c] = 8'hD0;
    buff [16'h04_2d] = 8'hE0;
    buff [16'h04_2e] = 8'hFA;
    buff [16'h04_2f] = 8'hD0;
    buff [16'h04_30] = 8'hE0;
    buff [16'h04_31] = 8'hF9;
    buff [16'h04_32] = 8'hD0;
    buff [16'h04_33] = 8'hE0;
    buff [16'h04_34] = 8'hF8;
    buff [16'h04_35] = 8'h12;
    buff [16'h04_36] = 8'h00;
    buff [16'h04_37] = 8'h89;
    buff [16'h04_38] = 8'hED;
    buff [16'h04_39] = 8'h64;
    buff [16'h04_3a] = 8'h80;
    buff [16'h04_3b] = 8'hFD;
    buff [16'h04_3c] = 8'h30;
    buff [16'h04_3d] = 8'hE7;
    buff [16'h04_3e] = 8'h01;
    buff [16'h04_3f] = 8'h1C;
    buff [16'h04_40] = 8'hD5;
    buff [16'h04_41] = 8'h83;
    buff [16'h04_42] = 8'hCB;
    buff [16'h04_43] = 8'hED;
    buff [16'h04_44] = 8'h33;
    buff [16'h04_45] = 8'hCC;
    buff [16'h04_46] = 8'h33;
    buff [16'h04_47] = 8'hF8;
    buff [16'h04_48] = 8'hD0;
    buff [16'h04_49] = 8'hE0;
    buff [16'h04_4a] = 8'hA2;
    buff [16'h04_4b] = 8'hE7;
    buff [16'h04_4c] = 8'h13;
    buff [16'h04_4d] = 8'h28;
    buff [16'h04_4e] = 8'hC3;
    buff [16'h04_4f] = 8'h13;
    buff [16'h04_50] = 8'hCC;
    buff [16'h04_51] = 8'h13;
    buff [16'h04_52] = 8'hFD;
    buff [16'h04_53] = 8'h22;
    buff [16'h04_54] = 8'h78;
    buff [16'h04_55] = 8'h7F;
    buff [16'h04_56] = 8'hE4;
    buff [16'h04_57] = 8'hF6;
    buff [16'h04_58] = 8'hD8;
    buff [16'h04_59] = 8'hFD;
    buff [16'h04_5a] = 8'h75;
    buff [16'h04_5b] = 8'h81;
    buff [16'h04_5c] = 8'h1B;
    buff [16'h04_5d] = 8'h02;
    buff [16'h04_5e] = 8'h00;
    buff [16'h04_5f] = 8'h03;
end

always @(posedge clk)
begin
  data1 <= #1 buff [addr];
  data2 <= #1 buff [addr+1];
  data3 <= #1 buff [addr+2];
end

endmodule
